
`include "inc.svh"

module top;

    initial begin
        `MY_DISPLAY ("Hello World!");
        $finish;
    end

endmodule

