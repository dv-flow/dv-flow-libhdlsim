module top;
    initial begin
        $display("VPI Test Start");
        #10;
        $display("VPI Test End");
        $finish;
    end
endmodule
