
module mod1_top;
    mod1 mod1_inst();

    initial begin
        $display("Hello World!");
    end

endmodule
