
`define MY_DISPLAY $display